//-- Fichero setbit.v
module setbit(output salida);
wire salida;

assign salida = 1;

endmodule
